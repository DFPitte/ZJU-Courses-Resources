`ifdef VERILATE
    localparam FILE_PATH = "initial.hex";
`else
    localparam FILE_PATH = "D:\\ZJU\\System\\sys1-sp24\\repo\\sys-project\\lab3-3\\syn\\initial.hex";//your initial.hex
`endif